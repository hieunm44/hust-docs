`timescale 1ns / 1ns

module main_tb;
	reg clk;
	// x: Phan thuc
	// y: Phan ao
	reg signed [15:0] xin [0:63];
	reg signed [15:0] yin [0:63];
	wire signed [15:0] xout [0:63];
	wire signed [15:0] yout [0:63];
	
	// Unit Under Test (UUT)
	main_cordic_fft uut (
		.clk(clk),
		
		.xin0(xin[0]), 
		.xin1(xin[1]), 
		.xin2(xin[2]), 
		.xin3(xin[3]), 
		.xin4(xin[4]), 
		.xin5(xin[5]),
		.xin6(xin[6]), 
		.xin7(xin[7]), 
		.xin8(xin[8]), 
		.xin9(xin[9]), 
		.xin10(xin[10]), 
		.xin11(xin[11]), 
		.xin12(xin[12]), 
		.xin13(xin[13]), 
		.xin14(xin[14]), 
		.xin15(xin[15]),
		.xin16(xin[16]), 
		.xin17(xin[17]), 
		.xin18(xin[18]), 
		.xin19(xin[19]), 
		.xin20(xin[20]), 
		.xin21(xin[21]), 
		.xin22(xin[22]), 
		.xin23(xin[23]), 
		.xin24(xin[24]), 
		.xin25(xin[25]), 
		.xin26(xin[26]), 
		.xin27(xin[27]), 
		.xin28(xin[28]), 
		.xin29(xin[29]), 
		.xin30(xin[30]), 
		.xin31(xin[31]), 
		.xin32(xin[32]), 
		.xin33(xin[33]), 
		.xin34(xin[34]), 
		.xin35(xin[35]), 
		.xin36(xin[36]), 
		.xin37(xin[37]), 
		.xin38(xin[38]), 
		.xin39(xin[39]), 
		.xin40(xin[40]), 
		.xin41(xin[41]), 
		.xin42(xin[42]), 
		.xin43(xin[43]), 
		.xin44(xin[44]), 
		.xin45(xin[45]), 
		.xin46(xin[46]), 
		.xin47(xin[47]), 
		.xin48(xin[48]), 
		.xin49(xin[49]), 
		.xin50(xin[50]), 
		.xin51(xin[51]), 
		.xin52(xin[52]), 
		.xin53(xin[53]), 
		.xin54(xin[54]), 
		.xin55(xin[55]), 
		.xin56(xin[56]), 
		.xin57(xin[57]), 
		.xin58(xin[58]), 
		.xin59(xin[59]), 
		.xin60(xin[60]), 
		.xin61(xin[61]), 
		.xin62(xin[62]), 
		.xin63(xin[63]), 
		
		.yin0(yin[0]), 
		.yin1(yin[1]), 
		.yin2(yin[2]), 
		.yin3(yin[3]), 
		.yin4(yin[4]), 
		.yin5(yin[5]),
		.yin6(yin[6]), 
		.yin7(yin[7]), 
		.yin8(yin[8]), 
		.yin9(yin[9]), 
		.yin10(yin[10]), 
		.yin11(yin[11]), 
		.yin12(yin[12]), 
		.yin13(yin[13]), 
		.yin14(yin[14]), 
		.yin15(yin[15]),
		.yin16(yin[16]), 
		.yin17(yin[17]), 
		.yin18(yin[18]), 
		.yin19(yin[19]), 
		.yin20(yin[20]), 
		.yin21(yin[21]), 
		.yin22(yin[22]), 
		.yin23(yin[23]), 
		.yin24(yin[24]), 
		.yin25(yin[25]), 
		.yin26(yin[26]), 
		.yin27(yin[27]), 
		.yin28(yin[28]), 
		.yin29(yin[29]), 
		.yin30(yin[30]), 
		.yin31(yin[31]), 
		.yin32(yin[32]), 
		.yin33(yin[33]), 
		.yin34(yin[34]), 
		.yin35(yin[35]), 
		.yin36(yin[36]), 
		.yin37(yin[37]), 
		.yin38(yin[38]), 
		.yin39(yin[39]), 
		.yin40(yin[40]), 
		.yin41(yin[41]), 
		.yin42(yin[42]), 
		.yin43(yin[43]), 
		.yin44(yin[44]), 
		.yin45(yin[45]), 
		.yin46(yin[46]), 
		.yin47(yin[47]), 
		.yin48(yin[48]), 
		.yin49(yin[49]), 
		.yin50(yin[50]), 
		.yin51(yin[51]), 
		.yin52(yin[52]), 
		.yin53(yin[53]), 
		.yin54(yin[54]), 
		.yin55(yin[55]), 
		.yin56(yin[56]), 
		.yin57(yin[57]), 
		.yin58(yin[58]), 
		.yin59(yin[59]), 
		.yin60(yin[60]), 
		.yin61(yin[61]), 
		.yin62(yin[62]), 
		.yin63(yin[63]), 
		
		.xout0(xout[0]), 
		.xout1(xout[1]), 
		.xout2(xout[2]), 
		.xout3(xout[3]), 
		.xout4(xout[4]), 
		.xout5(xout[5]),
		.xout6(xout[6]), 
		.xout7(xout[7]), 
		.xout8(xout[8]), 
		.xout9(xout[9]), 
		.xout10(xout[10]), 
		.xout11(xout[11]), 
		.xout12(xout[12]), 
		.xout13(xout[13]), 
		.xout14(xout[14]), 
		.xout15(xout[15]),
		.xout16(xout[16]), 
		.xout17(xout[17]), 
		.xout18(xout[18]), 
		.xout19(xout[19]), 
		.xout20(xout[20]), 
		.xout21(xout[21]), 
		.xout22(xout[22]), 
		.xout23(xout[23]), 
		.xout24(xout[24]), 
		.xout25(xout[25]), 
		.xout26(xout[26]), 
		.xout27(xout[27]), 
		.xout28(xout[28]), 
		.xout29(xout[29]), 
		.xout30(xout[30]), 
		.xout31(xout[31]), 
		.xout32(xout[32]), 
		.xout33(xout[33]), 
		.xout34(xout[34]), 
		.xout35(xout[35]), 
		.xout36(xout[36]), 
		.xout37(xout[37]), 
		.xout38(xout[38]), 
		.xout39(xout[39]), 
		.xout40(xout[40]), 
		.xout41(xout[41]), 
		.xout42(xout[42]), 
		.xout43(xout[43]), 
		.xout44(xout[44]), 
		.xout45(xout[45]), 
		.xout46(xout[46]), 
		.xout47(xout[47]), 
		.xout48(xout[48]), 
		.xout49(xout[49]), 
		.xout50(xout[50]), 
		.xout51(xout[51]), 
		.xout52(xout[52]), 
		.xout53(xout[53]), 
		.xout54(xout[54]), 
		.xout55(xout[55]), 
		.xout56(xout[56]), 
		.xout57(xout[57]), 
		.xout58(xout[58]), 
		.xout59(xout[59]), 
		.xout60(xout[60]), 
		.xout61(xout[61]), 
		.xout62(xout[62]), 
		.xout63(xout[63]), 
		
		.yout0(yout[0]), 
		.yout1(yout[1]), 
		.yout2(yout[2]), 
		.yout3(yout[3]), 
		.yout4(yout[4]), 
		.yout5(yout[5]),
		.yout6(yout[6]), 
		.yout7(yout[7]), 
		.yout8(yout[8]), 
		.yout9(yout[9]), 
		.yout10(yout[10]), 
		.yout11(yout[11]), 
		.yout12(yout[12]), 
		.yout13(yout[13]), 
		.yout14(yout[14]), 
		.yout15(yout[15]),
		.yout16(yout[16]), 
		.yout17(yout[17]), 
		.yout18(yout[18]), 
		.yout19(yout[19]), 
		.yout20(yout[20]), 
		.yout21(yout[21]), 
		.yout22(yout[22]), 
		.yout23(yout[23]), 
		.yout24(yout[24]), 
		.yout25(yout[25]), 
		.yout26(yout[26]), 
		.yout27(yout[27]), 
		.yout28(yout[28]), 
		.yout29(yout[29]), 
		.yout30(yout[30]), 
		.yout31(yout[31]), 
		.yout32(yout[32]), 
		.yout33(yout[33]), 
		.yout34(yout[34]), 
		.yout35(yout[35]), 
		.yout36(yout[36]), 
		.yout37(yout[37]), 
		.yout38(yout[38]), 
		.yout39(yout[39]), 
		.yout40(yout[40]), 
		.yout41(yout[41]), 
		.yout42(yout[42]), 
		.yout43(yout[43]), 
		.yout44(yout[44]), 
		.yout45(yout[45]), 
		.yout46(yout[46]), 
		.yout47(yout[47]), 
		.yout48(yout[48]), 
		.yout49(yout[49]), 
		.yout50(yout[50]), 
		.yout51(yout[51]), 
		.yout52(yout[52]), 
		.yout53(yout[53]), 
		.yout54(yout[54]), 
		.yout55(yout[55]), 
		.yout56(yout[56]), 
		.yout57(yout[57]), 
		.yout58(yout[58]), 
		.yout59(yout[59]), 
		.yout60(yout[60]), 
		.yout61(yout[61]), 
		.yout62(yout[62]), 
		.yout63(yout[63])
	);
	
	
	integer i;
	initial
	begin
		//Khoi tao cac dau vao =0
		for (i=0;i<64;i=i+1)
		begin
			xin[i]=0;
			yin[i]=0;
		end
	
		#100;        
		// Thiet lap cac gia tri dau vao
		
		xin[0]=1000;
		xin[1]=-800;
		xin[2]=1000;
		xin[3]=-800;
		xin[4]=1000;
		xin[5]=-800;
		xin[6]=1000;
		xin[7]=-800;
		xin[8]=1000;
		xin[9]=-800;
		xin[10]=1000;
		xin[11]=-800;
		xin[12]=1000;
		xin[13]=-800;
		xin[14]=1000;
		xin[15]=-800;
		xin[16]=1000;
		xin[17]=-800;
		xin[18]=1000;
		xin[19]=-800;
		xin[20]=1000;
		xin[21]=-800;
		xin[22]=1000;
		xin[23]=-800;
		xin[24]=1000;
		xin[25]=-800;
		xin[26]=1000;
		xin[27]=-800;
		xin[28]=1000;
		xin[29]=-800;
		xin[30]=1000;
		xin[31]=-800;
		/*
		xin[32]=420;
		xin[33]=430;
		xin[34]=440;
		xin[35]=450;
		xin[36]=460;
		xin[37]=470;
		xin[38]=480;
		xin[39]=490;
		xin[40]=500;
		xin[41]=510;
		xin[42]=520;
		xin[43]=530;
		xin[44]=540;
		xin[45]=550;
		xin[46]=560;
		xin[47]=570;
		xin[48]=580;
		xin[49]=590;
		xin[50]=600;
		xin[51]=610;
		xin[52]=620;
		xin[53]=630;
		xin[54]=640;
		xin[55]=650;
		xin[56]=660;
		xin[57]=670;
		xin[58]=680;
		xin[59]=690;
		xin[60]=700;
		xin[61]=710;
		xin[62]=720;
		xin[63]=730;
		
		/*
		xin[0]=3200;
		xin[1]=3200;
		xin[2]=3200;
		xin[3]=3200;
		xin[4]=3200;
		xin[5]=3200;
		xin[6]=3200;
		xin[7]=3200;
		*/
		
		yin[0]=0;
		yin[1]=0;
		yin[2]=0;
		yin[3]=0;
		yin[4]=0;
		yin[5]=0;
		yin[6]=0;
		yin[7]=0;
		yin[8]=0;
		yin[9]=0;
		yin[10]=0;
		yin[11]=0;
		yin[12]=0;
		yin[13]=0;
		yin[14]=0;
		yin[15]=0;
		yin[16]=0;
		yin[17]=0;
		yin[18]=0;
		yin[19]=0;
		yin[20]=0;
		yin[21]=0;
		yin[22]=0;
		yin[23]=0;
		yin[24]=0;
		yin[25]=0;
		yin[26]=0;
		yin[27]=0;
		yin[28]=0;
		yin[29]=0;
		yin[30]=0;
		yin[31]=0;
		yin[32]=0;
		yin[33]=0;
		yin[34]=0;
		yin[35]=0;
		yin[36]=0;
		yin[37]=0;
		yin[38]=0;
		yin[39]=0;
		yin[40]=0;
		yin[41]=0;
		yin[42]=0;
		yin[43]=0;
		yin[44]=0;
		yin[45]=0;
		yin[46]=0;
		yin[47]=0;
		yin[48]=0;
		yin[49]=0;
		yin[50]=0;
		yin[51]=0;
		yin[52]=0;
		yin[53]=0;
		yin[54]=0;
		yin[55]=0;
		yin[56]=0;
		yin[57]=0;
		yin[58]=0;
		yin[59]=0;
		yin[60]=0;
		yin[61]=0;
		yin[62]=0;
		yin[63]=0;

		#1000;
		
		// Hien thi ket qua tren Transcript
		$display("x[0]=%d %di\nx[1]=%d %di\nx[2]=%d %di\nx[3]=%d %di\nx[4]=%d %di\nx[5]=%d %di\nx[6]=%d %di\nx[7]=%d %di\nx[8]=%d %di\nx[9]=%d %di\nx[10]=%d %di\nx[11]=%d %di\nx[12]=%d %di\nx[13]=%d %di\nx[14]=%d %di\nx[15]=%d %di\nx[16]=%d %di\nx[17]=%d %di\nx[18]=%d %di\nx[19]=%d %di\nx[20]=%d %di\nx[21]=%d %di\nx[22]=%d %di\nx[23]=%d %di\nx[24]=%d %di\nx[25]=%d %di\nx[26]=%d %di\nx[27]=%d %di\nx[28]=%d %di\nx[29]=%d %di\nx[30]=%d %di\nx[31]=%d %di\nx[32]=%d %di\nx[33]=%d %di\nx[34]=%d %di\nx[35]=%d %di\nx[36]=%d %di\nx[37]=%d %di\nx[38]=%d %di\nx[39]=%d %di\nx[40]=%d %di\nx[41]=%d %di\nx[42]=%d %di\nx[43]=%d %di\nx[44]=%d %di\nx[45]=%d %di\nx[46]=%d %di\nx[47]=%d %di\nx[48]=%d %di\nx[49]=%d %di\nx[50]=%d %di\nx[51]=%d %di\nx[52]=%d %di\nx[53]=%d %di\nx[54]=%d %di\nx[55]=%d %di\nx[56]=%d %di\nx[57]=%d %di\nx[58]=%d %di\nx[59]=%d %di\nx[60]=%d %di\nx[61]=%d %di\nx[62]=%d %di\nx[63]=%d %di\n\n",xin[0],yin[0],xin[1],yin[1],xin[2],yin[2],xin[3],yin[3],xin[4],yin[4],xin[5],yin[5],xin[6],yin[6],xin[7],yin[7],xin[8],yin[8],xin[9],yin[9],xin[10],yin[10],xin[11],yin[11],xin[12],yin[12],xin[13],yin[13],xin[14],yin[14],xin[15],yin[15],xin[16],yin[16],xin[17],yin[17],xin[18],yin[18],xin[19],yin[19],xin[20],yin[20],xin[21],yin[21],xin[22],yin[22],xin[23],yin[23],xin[24],yin[24],xin[25],yin[25],xin[26],yin[26],xin[27],yin[27],xin[28],yin[28],xin[29],yin[29],xin[30],yin[30],xin[31],yin[31],xin[32],yin[32],xin[33],yin[33],xin[34],yin[34],xin[35],yin[35],xin[36],yin[36],xin[37],yin[37],xin[38],yin[38],xin[39],yin[39],xin[40],yin[40],xin[41],yin[41],xin[42],yin[42],xin[43],yin[43],xin[44],yin[44],xin[45],yin[45],xin[46],yin[46],xin[47],yin[47],xin[48],yin[48],xin[49],yin[49],xin[50],yin[50],xin[51],yin[51],xin[52],yin[52],xin[53],yin[53],xin[54],yin[54],xin[55],yin[55],xin[56],yin[56],xin[57],yin[57],xin[58],yin[58],xin[59],yin[59],xin[60],yin[60],xin[61],yin[61],xin[62],yin[62],xin[63],yin[63]);
		$display("X[0]=%d %di\nX[1]=%d %di\nX[2]=%d %di\nX[3]=%d %di\nX[4]=%d %di\nX[5]=%d %di\nX[6]=%d %di\nX[7]=%d %di\nX[8]=%d %di\nX[9]=%d %di\nX[10]=%d %di\nX[11]=%d %di\nX[12]=%d %di\nX[13]=%d %di\nX[14]=%d %di\nX[15]=%d %di\nX[16]=%d %di\nX[17]=%d %di\nX[18]=%d %di\nX[19]=%d %di\nX[20]=%d %di\nX[21]=%d %di\nX[22]=%d %di\nX[23]=%d %di\nX[24]=%d %di\nX[25]=%d %di\nX[26]=%d %di\nX[27]=%d %di\nX[28]=%d %di\nX[29]=%d %di\nX[30]=%d %di\nX[31]=%d %di\nX[32]=%d %di\nX[33]=%d %di\nX[34]=%d %di\nX[35]=%d %di\nX[36]=%d %di\nX[37]=%d %di\nX[38]=%d %di\nX[39]=%d %di\nX[40]=%d %di\nX[41]=%d %di\nX[42]=%d %di\nX[43]=%d %di\nX[44]=%d %di\nX[45]=%d %di\nX[46]=%d %di\nX[47]=%d %di\nX[48]=%d %di\nX[49]=%d %di\nX[50]=%d %di\nX[51]=%d %di\nX[52]=%d %di\nX[53]=%d %di\nX[54]=%d %di\nX[55]=%d %di\nX[56]=%d %di\nX[57]=%d %di\nX[58]=%d %di\nX[59]=%d %di\nX[60]=%d %di\nX[61]=%d %di\nX[62]=%d %di\nX[63]=%d %di\n\n",xout[0],yout[0],xout[1],yout[1],xout[2],yout[2],xout[3],yout[3],xout[4],yout[4],xout[5],yout[5],xout[6],yout[6],xout[7],yout[7],xout[8],yout[8],xout[9],yout[9],xout[10],yout[10],xout[11],yout[11],xout[12],yout[12],xout[13],yout[13],xout[14],yout[14],xout[15],yout[15],xout[16],yout[16],xout[17],yout[17],xout[18],yout[18],xout[19],yout[19],xout[20],yout[20],xout[21],yout[21],xout[22],yout[22],xout[23],yout[23],xout[24],yout[24],xout[25],yout[25],xout[26],yout[26],xout[27],yout[27],xout[28],yout[28],xout[29],yout[29],xout[30],yout[30],xout[31],yout[31],xout[32],yout[32],xout[33],yout[33],xout[34],yout[34],xout[35],yout[35],xout[36],yout[36],xout[37],yout[37],xout[38],yout[38],xout[39],yout[39],xout[40],yout[40],xout[41],yout[41],xout[42],yout[42],xout[43],yout[43],xout[44],yout[44],xout[45],yout[45],xout[46],yout[46],xout[47],yout[47],xout[48],yout[48],xout[49],yout[49],xout[50],yout[50],xout[51],yout[51],xout[52],yout[52],xout[53],yout[53],xout[54],yout[54],xout[55],yout[55],xout[56],yout[56],xout[57],yout[57],xout[58],yout[58],xout[59],yout[59],xout[60],yout[60],xout[61],yout[61],xout[62],yout[62],xout[63],yout[63]);
	end
	
	// Thiet lap xung clock
	initial
	begin
		clk=1'b0;
		forever #5 clk=~clk;
	end
    

endmodule