CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 75 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 171 457 268
110100498 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 218 261 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4212 0 0
2
42074.7 1
0
13 Logic Switch~
5 218 216 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4720 0 0
2
42074.7 0
0
13 Logic Switch~
5 217 171 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5551 0 0
2
42074.7 0
0
9 2-In AND~
219 716 216 0 3 22
0 4 3 2
0
0 0 368 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6986 0 0
2
42074.7 0
0
9 2-In AND~
219 485 251 0 3 22
0 8 7 6
0
0 0 368 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
8745 0 0
2
42074.7 0
0
9 2-In AND~
219 482 178 0 3 22
0 8 10 5
0
0 0 368 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9592 0 0
2
42074.7 0
0
8 2-In OR~
219 599 189 0 3 22
0 5 9 4
0
0 0 368 0
6 74LS32
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8748 0 0
2
42074.7 0
0
9 Inverter~
13 352 215 0 2 22
0 11 9
0
0 0 368 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 1 0
1 U
7168 0 0
2
42074.7 0
0
14 Logic Display~
6 775 140 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
631 0 0
2
42074.7 0
0
9 Inverter~
13 354 259 0 2 22
0 10 7
0
0 0 368 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 1 0
1 U
9466 0 0
2
42074.7 0
0
8 2-In OR~
219 599 245 0 3 22
0 9 6 3
0
0 0 368 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3266 0 0
2
42074.7 0
0
9 Inverter~
13 351 171 0 2 22
0 12 8
0
0 0 368 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 250
65 0 0 0 6 1 1 0
1 U
7693 0 0
2
42074.7 0
0
14
3 1 2 0 0 8320 0 4 9 0 0 3
737 216
775 216
775 158
3 2 3 0 0 4224 0 11 4 0 0 4
632 245
684 245
684 225
692 225
1 3 4 0 0 4224 0 4 7 0 0 4
692 207
640 207
640 189
632 189
3 1 5 0 0 4224 0 6 7 0 0 4
503 178
578 178
578 180
586 180
3 2 6 0 0 4224 0 5 11 0 0 4
506 251
578 251
578 254
586 254
2 2 7 0 0 4224 0 10 5 0 0 4
375 259
440 259
440 260
461 260
0 1 8 0 0 4224 0 0 5 13 0 3
406 171
406 242
461 242
1 0 9 0 0 8192 0 11 0 0 9 3
586 236
577 236
577 215
2 2 9 0 0 4224 0 8 7 0 0 4
373 215
578 215
578 198
586 198
0 2 10 0 0 8320 0 0 6 11 0 5
262 261
262 186
438 186
438 187
458 187
1 1 10 0 0 0 0 1 10 0 0 4
230 261
331 261
331 259
339 259
1 1 11 0 0 4224 0 2 8 0 0 4
230 216
329 216
329 215
337 215
2 1 8 0 0 0 0 12 6 0 0 4
372 171
443 171
443 169
458 169
1 1 12 0 0 4224 0 3 12 0 0 2
229 171
336 171
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
151 246 180 270
157 250 173 266
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
147 208 176 232
153 212 169 228
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
144 158 173 182
150 162 166 178
2 S1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
