CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 75 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
176 411 1364 747
110100498 0
0
6 Title:
5 Name:
0
0
0
5
6 74LS90
107 510 231 0 10 21
0 2 2 7 6 4 5 8 6 7
5
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 512 0 0 0 0
1 U
34 0 0
2
42074.8 0
0
14 Logic Display~
6 640 157 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
42074.8 0
0
7 Ground~
168 425 299 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8402 0 0
2
42074.8 0
0
14 Logic Display~
6 340 159 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3751 0 0
2
42074.8 0
0
7 Pulser~
4 259 260 0 10 12
0 9 10 3 4 0 0 10 10 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4292 0 0
2
42074.8 0
0
8
3 1 3 0 0 8320 0 5 4 0 0 3
283 251
340 251
340 177
4 5 4 0 0 4224 0 5 1 0 0 4
289 260
459 260
459 249
472 249
6 10 5 0 0 12416 0 1 1 0 0 6
472 258
463 258
463 278
555 278
555 258
542 258
1 0 6 0 0 8320 0 2 0 0 5 3
640 175
640 222
550 222
4 8 6 0 0 0 0 1 1 0 0 6
478 231
463 231
463 184
550 184
550 222
542 222
3 9 7 0 0 12416 0 1 1 0 0 6
478 222
468 222
468 273
550 273
550 240
542 240
2 0 2 0 0 4096 0 1 0 0 8 2
478 213
425 213
1 1 2 0 0 4224 0 3 1 0 0 3
425 293
425 204
478 204
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
