CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 75 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 171 457 268
110100498 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 412 110 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9442 0 0
2
42074.8 0
0
7 Ground~
168 422 251 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9424 0 0
2
42074.8 0
0
12 Hex Display~
7 699 189 0 18 19
10 6 7 8 9 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9968 0 0
2
42074.8 0
0
2 +V
167 620 121 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9281 0 0
2
42074.8 0
0
7 74LS168
8 526 242 0 14 29
0 2 2 3 10 11 12 13 5 4
14 9 8 7 6
0
0 0 4848 0
8 74LS168A
-28 -60 28 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 6 5 4 3 9 1
15 11 12 13 14 7 10 2 6 5
4 3 9 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
8464 0 0
2
42074.8 0
0
14 Logic Display~
6 339 164 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
42074.8 0
0
7 Pulser~
4 259 227 0 10 12
0 15 16 17 3 0 0 10 10 9
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3171 0 0
2
42074.8 0
0
10
1 0 3 0 0 4096 0 6 0 0 3 2
339 182
339 224
1 0 2 0 0 8320 0 2 0 0 4 3
422 245
422 210
488 210
3 4 3 0 0 4224 0 5 7 0 0 4
494 224
297 224
297 227
289 227
1 2 2 0 0 0 0 5 5 0 0 2
488 206
488 215
9 1 4 0 0 12416 0 5 1 0 0 4
558 215
568 215
568 110
424 110
8 1 5 0 0 8320 0 5 4 0 0 3
564 206
620 206
620 130
14 1 6 0 0 4224 0 5 3 0 0 3
558 278
708 278
708 213
13 2 7 0 0 4224 0 5 3 0 0 3
558 269
702 269
702 213
12 3 8 0 0 4224 0 5 3 0 0 3
558 260
696 260
696 213
11 4 9 0 0 4224 0 5 3 0 0 3
558 251
690 251
690 213
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
