CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 75 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 171 457 268
110100498 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 220 262 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
42074.8 0
0
13 Logic Switch~
5 218 216 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
5.89699e-315 0
0
13 Logic Switch~
5 217 171 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.89699e-315 0
0
7 Ground~
168 340 331 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3670 0 0
2
42074.8 0
0
2 +V
167 259 303 0 1 3
0 11
0
0 0 54256 90
2 5V
-8 -15 6 -7
2 V4
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5616 0 0
2
42074.8 0
0
7 74LS138
19 423 234 0 14 29
0 14 13 12 11 2 2 10 9 8
7 6 5 4 3
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
9323 0 0
2
42074.8 0
0
14 Logic Display~
6 799 76 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
42074.8 1
0
14 Logic Display~
6 754 80 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
42074.8 0
0
14 Logic Display~
6 714 82 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
42074.8 2
0
14 Logic Display~
6 666 89 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
42074.8 1
0
14 Logic Display~
6 628 86 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
42074.8 0
0
14 Logic Display~
6 597 95 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
42074.8 2
0
14 Logic Display~
6 562 91 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
42074.8 1
0
14 Logic Display~
6 534 86 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
42074.8 0
0
14 Logic Display~
6 338 93 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
42074.8 0
0
14 Logic Display~
6 305 94 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
42074.8 0
0
14 Logic Display~
6 267 96 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89699e-315 0
0
17
14 1 3 0 0 4224 0 6 7 0 0 3
461 270
799 270
799 94
1 13 4 0 0 8320 0 8 6 0 0 3
754 98
754 261
461 261
12 1 5 0 0 4224 0 6 9 0 0 3
461 252
714 252
714 100
1 11 6 0 0 8320 0 10 6 0 0 3
666 107
666 243
461 243
10 1 7 0 0 4224 0 6 11 0 0 3
461 234
628 234
628 104
9 1 8 0 0 4224 0 6 12 0 0 3
461 225
597 225
597 113
1 8 9 0 0 4224 0 13 6 0 0 3
562 109
562 216
461 216
7 1 10 0 0 8320 0 6 14 0 0 3
461 207
534 207
534 104
1 6 2 0 0 4224 0 4 6 0 0 3
340 325
340 270
385 270
6 5 2 0 0 0 0 6 6 0 0 2
385 270
385 261
4 1 11 0 0 4224 0 6 5 0 0 4
391 252
278 252
278 301
270 301
1 0 12 0 0 4224 0 15 0 0 15 2
338 111
338 262
1 0 13 0 0 4096 0 16 0 0 16 4
305 112
305 211
306 211
306 216
1 0 14 0 0 4096 0 17 0 0 17 2
267 114
267 171
1 3 12 0 0 0 0 1 6 0 0 4
232 262
356 262
356 225
391 225
1 2 13 0 0 4224 0 2 6 0 0 2
230 216
391 216
1 1 14 0 0 4224 0 3 6 0 0 4
229 171
361 171
361 207
391 207
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
151 244 180 268
157 248 173 264
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
144 158 173 182
150 162 166 178
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
147 208 176 232
153 212 169 228
2 S2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
